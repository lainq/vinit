module utility

pub fn helloworld() {
	println("Hello")
}