module argparse
