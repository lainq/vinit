module main

pub fn helloworld() {
	println("Hello")
}