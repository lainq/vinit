module vinit
